library ieee;
use ieee.std_logic_1164.all;

package cte_tipos_UF_pkg is 

-- ALU OPCODES
constant ALU_MOVI: std_logic := '0';
constant ALU_MOVHI: std_logic := '1';
-- --
       
constant PE:  std_logic:= '1';

END PACKAGE cte_tipos_UF_pkg;